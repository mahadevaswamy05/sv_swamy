 Hi ,
