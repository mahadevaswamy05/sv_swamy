10000
10001
10010


This is Mahadevaswamy
from Bengalore
