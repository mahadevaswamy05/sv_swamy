This is Mahadevaswamy
from Bengalore
